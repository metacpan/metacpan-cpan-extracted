Animal|Vegetable\|Mineral|Description
