Minst net1
+ net2 net3
+ net4 nmos l=0.09u
+ w=0.13u
.END

*This line is not read
