
module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule


module my_mod ( port1 , port2 , port3, porta, portb, portc
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, port_yada , port_bingo , port_bango , port_x , port_y , port_z
	, port1abcd , porsdfdt2 , portfdfsdf3, portasdfdf, portbadfd, portcsdf
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
	, \m_esc_nameaa!3!332 , \m_esc_namebb!3!33 , \m_esc_namecc!3!323 
 
 );

   mod_name inst_name ( 
	  .port({n111, n222, n333, n444, n555, n666 , n777, n888})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	, .yet_another_port({a_big_port, some_big_port, a_port, b_port, c_port
	, port_yada, \mport_bin!2!45go, port_bango, \mport_dod1!3!o, port_of_call})
	);

endmodule

