Animal|Vegetable\|Mineral|Description
Wombat|Celery or asparagus|Cute and\nfurry
Moose|Choco\late|C:\\Delicious
