Animal|Vegetable\|Mineral|Description
Wombat|Celery or asparagus|Cute and\nfurry
Moose|Chocolate|C:\\Delicious
